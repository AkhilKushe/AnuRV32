module sigExt ( data_in,
		data_out);

parameter WIDTH = 8;
input [WIDTH-1:0] data_in;
output [31:0] data_out;

//Sign extend data_in to 32 bits
assign data_out = {{(32-WIDTH){data_in[WIDTH-1]}} , data_in};

endmodule

module zeroExt ( data_in,
		data_out);
parameter WIDTH = 8;
input [WIDTH -1 : 0] data_in;
output [31:0] data_out;

//Zero extend data_in to 32 bits
assign data_out = {{(32-WIDTH){1'b0}} , data_in};

endmodule

module extend32 ( data_in,
		sig,
		b_hbar,
		bypass,
		data_out);

input [31:0] data_in;
input sig, b_hbar, bypass;
output reg [31:0] data_out;

wire [31:0] z_extend8_w;
wire [31:0] z_extend16_w;
wire [31:0] s_extend8_w;
wire [31:0] s_extend16_w;

zeroExt #(.WIDTH(8)) zE8(.data_in(data_in[7:0]), .data_out(z_extend8_w));
zeroExt #(.WIDTH(16)) zE16(.data_in(data_in[15:0]), .data_out(z_extend16_w));
sigExt #(.WIDTH(8)) sE8(.data_in(data_in[7:0]), .data_out(s_extend8_w));
sigExt #(.WIDTH(16)) sE16(.data_in(data_in[15:0]), .data_out(s_extend16_w));

always @(*) begin
	if (bypass) begin
		data_out = data_in;
	end else begin
		if (b_hbar) begin
			if (sig) begin
				data_out = s_extend8_w;
			end else begin
				data_out = z_extend8_w;
			end
		end else begin
			if (sig) begin
				data_out = s_extend16_w;
			end else begin
				data_out = z_extend16_w;
			end
		end
	end

end

endmodule

