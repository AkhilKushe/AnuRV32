package agent_pkg; 
    import uvm_pkg::*; 
    `include "monitor.sv"
    `include "agent.sv"
endpackage